`timescale 1ns / 1ps

module tb_ripple_carry_adder_32bit;
    reg [31:0] a, b;
    reg c_in;
    wire [31:0] sum;
    wire c_out;
    
    ripple_carry_adder_src dut(.a(a),.b(b),.c_in(c_in),.sum(sum),.c_out(c_out));
    
    initial begin
        a = 32'b00000000000000000000000000000000;
        b = 32'b00000000000000000000000000000000;
        c_in = 0;
        
        #20
        a = 32'b11110111001010111110010101001111;
        b = 32'b10010111100101011111000110010101;
        c_in = 1;

        #20
        a = 32'b01001110100101001111101001011100;
        b = 32'b11001011010011001110101000110100;
        c_in = 0;

        #20
        a = 32'b01111010111001011001101111011011;
        b = 32'b00101101001001010101011000110101;
        c_in = 1;

        #20
        a = 32'b10101010001011011001111001101110;
        b = 32'b11011111111100000101010111011101;
        c_in = 0;

        #20
        a = 32'b10101001101101101101101101000101;
        b = 32'b10110001101101011100111000101111;
        c_in = 1;

        #20
        a = 32'b11101110111011001100110110101001;
        b = 32'b11111001001100110001111011101111;
        c_in = 0;

        #20
        a = 32'b01110000111001011011010010011110;
        b = 32'b01101011011011011011010110010110;
        c_in = 1;

        #20
        a = 32'b10101010111011101010001101001100;
        b = 32'b11110110010001101110011001100101;
        c_in = 0;

        #20
        a = 32'b11101111010011110110100101001010;
        b = 32'b01101011010000110010110111001110;
        c_in = 1;

        #20
        a = 32'b10101100111010001001001001010100;
        b = 32'b11101011001011001100111000111000;
        c_in = 0;

        #20
        a = 32'b11100110100111110011100111000101;
        b = 32'b11011101010000111010111110010010;
        c_in = 1;

        #20
        a = 32'b11001111011010111110101110111100;
        b = 32'b01011111110111010110010111011000;
        c_in = 0;

        #20
        a = 32'b01001011101010001010110110001000;
        b = 32'b11010010101101110011110001001011;
        c_in = 1;

        #20
        a = 32'b11101000111011011001110110110111;
        b = 32'b10001001111100101111000101101010;
        c_in = 0;

        #20
        a = 32'b11011111110010101100100101001110;
        b = 32'b10010010101010101010111111010101;
        c_in = 1;
        
        #20 $finish;
    end
endmodule
