// TODO: change these paths if you move the Memory or RegFile instantiation
// to a different module
`define RF_PATH   CPU.icpu.rf
`define DMEM_PATH CPU.imem
`define IMEM_PATH CPU.imem
